
module audio_controller (
    input wire clk,
    input wire rst,
    input wire [2:0] button_press,
    output wire AUD_XCK,
    output wire AUD_DACDAT,
    inout wire AUD_DACLRCK,
    inout wire AUD_BCLK,
    output wire FPGA_I2C_SCLK,
    inout wire FPGA_I2C_SDAT
);

    // Audio frequencies for each column
    parameter FREQ_LEFT   = 500;   // A5 note
	 
    parameter FREQ_MIDDLE = 700;  // C6 note
	 
    parameter FREQ_RIGHT  = 900;  // D6 note

    // Clock generation
    wire audio_clk;   // 12.288 MHz clock for WM8731
	 
    wire sample_clk;  // Audio sample clock
	 

    // Audio data signals
    reg [15:0] audio_data;
	 
    reg data_valid;

    // Sine wave phase accumulators
    reg [31:0] phase_accum_left;
	 
    reg [31:0] phase_accum_middle;
	 
    reg [31:0] phase_accum_right;

    // Frequency increment calculations
    wire [31:0] freq_inc_left   = 32'h100000 * FREQ_LEFT / 48000;
	 
    wire [31:0] freq_inc_middle = 32'h100000 * FREQ_MIDDLE / 48000;
	 
    wire [31:0] freq_inc_right  = 32'h100000 * FREQ_RIGHT / 48000;

    // Audio PLL and codec configuration modules
    audio_pll pll_inst (
        .inclk0(clk),
        .c0(audio_clk),
        .c1(sample_clk)
    );

    codec_config codec_config_inst (
        .clk(clk),
        .rst(rst),
        .FPGA_I2C_SCLK(FPGA_I2C_SCLK),
        .FPGA_I2C_SDAT(FPGA_I2C_SDAT)
    );

    // Audio data generation
    always @(posedge sample_clk or posedge rst) begin
        if (rst) begin
            phase_accum_left <= 0;
            phase_accum_middle <= 0;
            phase_accum_right <= 0;
            audio_data <= 16'd0;
            data_valid <= 1'b0;
        end else begin
            // Update phase accumulators when buttons are pressed
            if (button_press[0]) begin
                phase_accum_left <= phase_accum_left + freq_inc_left;
            end else begin
                phase_accum_left <= 0;
            end

            if (button_press[1]) begin
                phase_accum_middle <= phase_accum_middle + freq_inc_middle;
            end else begin
                phase_accum_middle <= 0;
            end

            if (button_press[2]) begin
                phase_accum_right <= phase_accum_right + freq_inc_right;
            end else begin
                phase_accum_right <= 0;
            end

            // Mix audio outputs
            if (button_press != 3'b000) begin
                audio_data <= {
                    sine_lookup(phase_accum_left[31:24]),
                    sine_lookup(phase_accum_middle[31:24])
                };
                data_valid <= 1'b1;
            end else begin
                audio_data <= 16'd0;
                data_valid <= 1'b0;
            end
        end
    end

    // I2S transmitter
    i2s_transmitter i2s_tx_inst (
        .clk(audio_clk),
        .rst(rst),
        .data_in(audio_data),
        .data_valid(data_valid),
        .BCLK(AUD_BCLK),
        .LRCLK(AUD_DACLRCK),
        .DACDAT(AUD_DACDAT)
    );

    // Master clock generation for WM8731
    assign AUD_XCK = audio_clk;

    // Sine wave lookup function (8-bit resolution)
    function [7:0] sine_lookup;
        input [7:0] phase;
        begin
            case(phase[7:6])
                2'b00: sine_lookup = {1'b0, phase[6:0]} + 8'd128;       // 0 to π/2
                2'b01: sine_lookup = 8'd255 - {1'b0, phase[6:0]};       // π/2 to π
                2'b10: sine_lookup = ~{1'b0, phase[6:0]} + 8'd128;      // π to 3π/2
                2'b11: sine_lookup = {1'b0, phase[6:0]} + 8'd1;         // 3π/2 to 2π
            endcase
        end
    endfunction
endmodule

// I2S Transmitter Module
module i2s_transmitter (
    input wire clk,           // Audio bit clock
    input wire rst,           // Reset signal
    input wire [15:0] data_in,// Audio data to transmit
    input wire data_valid,    // Data valid flag
    
    inout wire BCLK,          // Bit clock
    inout wire LRCLK,         // Left/Right clock
    output reg DACDAT         // Serial audio data
);
    reg [4:0] bit_count;
    reg lr_select;

    // Bit clock generation (toggling)
    assign BCLK = clk;

    // Left/Right clock generation
    assign LRCLK = lr_select;

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            bit_count <= 5'd0;
            lr_select <= 1'b0;
            DACDAT <= 1'b0;
        end else begin
            // Left/Right clock toggles every 16 bits
            if (bit_count == 5'd0) begin
                lr_select <= ~lr_select;
            end

            // Transmit data when valid
            if (data_valid) begin
                if (bit_count < 5'd16) begin
                    DACDAT <= data_in[15 - bit_count];
                    bit_count <= bit_count + 1'b1;
                end else begin
                    bit_count <= 5'd0;
                end
            end else begin
                bit_count <= 5'd0;
                DACDAT <= 1'b0;
            end
        end
    end
endmodule

// Codec Configuration Module (Simplified)
module codec_config (
    input wire clk,
    input wire rst,
    output wire FPGA_I2C_SCLK,
    inout wire FPGA_I2C_SDAT
);
    // Placeholder for codec initialization 
    // In a real implementation, you'd send I2C configuration 
    // commands to set up the WM8731 codec
    assign FPGA_I2C_SCLK = 1'b1;
    assign FPGA_I2C_SDAT = 1'bz;
endmodule

// Audio PLL Module (Placeholder)
module audio_pll (
    input wire inclk0,
    output wire c0,  // 12.288 MHz for audio master clock
    output wire c1   // 48 kHz sample clock
);
    // For simulation, we'll use simple assignments
    assign c0 = inclk0;  // Simplified clock generation
    assign c1 = inclk0;  // Simplified sample clock
endmodule
